`timescale 1ns / 1ps

module forwarding_unit(
    input logic [4:0] id_ex_rs1, id_ex_rs2,
    input logic [4:0] ex_mem_rd,
    input logic [4:0] mem_wb_rd,
    input logic ex_mem_regwrite,
    input logic mem_wb_regwrite,
    output logic [1:0] forwardA,
    output logic [1:0] forwardB
);
    always_comb begin
        forwardA = 2'b00;
        forwardB = 2'b00;
        if (ex_mem_regwrite && (ex_mem_rd != 0)) begin
            if (ex_mem_rd == id_ex_rs1) forwardA = 2'b10;
            if (ex_mem_rd == id_ex_rs2) forwardB = 2'b10;
        end
        if (mem_wb_regwrite && (mem_wb_rd != 0)) begin
            if (!(ex_mem_regwrite && (ex_mem_rd != 0) && (ex_mem_rd == id_ex_rs1)) &&
                 (mem_wb_rd == id_ex_rs1)) forwardA = 2'b01;

            if (!(ex_mem_regwrite && (ex_mem_rd != 0) && (ex_mem_rd == id_ex_rs2)) &&
                 (mem_wb_rd == id_ex_rs2)) forwardB = 2'b01;
        end
    end

endmodule
